module or_gate ( input x1, x2, output out );
  
  assign
      out   = x1 | x2 ; 
    
endmodule