module or_gate_3 ( input x1, x2, x3, output  out );
  
  assign
      out   = x1 | x2 | x3 ; 
    
endmodule