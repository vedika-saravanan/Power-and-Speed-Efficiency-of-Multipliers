module or_gate_4 ( input x1, x2,x3, x4, output out );
  
  assign
      out   = x1 | x2 | x3 | x4 ; 
    
endmodule